`timescale 1ns / 1ns
 
module tb_horse_race_lamp;

    // Inputs
    reg [1:0] S;        // ??????
    reg clk;             // ????
    reg reset;           // ????

    // Outputs
    wire [7:0] Y;       // LED???

    // ?????????UUT?
    horse_race_lamp uut (
        .S(S),
        .clk(clk),
        .reset(reset),
        .Y(Y)
    );

    // ??????
    initial begin
        clk = 0;   // ??????0
        forever #5 clk = ~clk;  // ?5?????????
    end

    // ????????
    initial begin
        $display("Running testbench");

        // ?????
        reset = 1;  // ?????????
        S = 2'b00;   // ?????00
        #10 reset = 0;  // ????
        #400;         // ??400????

        // ???????
        reset = 1; 
        #5 reset = 0;  // ??????5????
        S = 2'b01;     // ?????01
        #200;          // ??200????

        reset = 1;
        #5 reset = 0;
        S = 2'b10;     // ?????10
        #200;          // ??200????

        reset = 1;
        #5 reset = 0;
        S = 2'b11;     // ?????11
        #100;          // ??100????

        $stop;         // ????
    end

endmodule
